--Square
library ieee;
use ieee.std_logic_1164.all;

entity SquareSquarer is
	Port(
		b:	in std_logic_vector(15 downto 0);
		y:	out std_logic_vector(31 downto 0)
		);
end SquareSquarer;

architecture Behavioral of SquareSquarer is

begin
y(23) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(22) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(21) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0));
y(20) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0)));
y(19) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0));
y(18) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0)));
y(17) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0)));
y(16) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(15) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0)));
y(14) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(13) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(12) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(11) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(10) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(9) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(8) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and (not b(0)));
y(7) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
y(6) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0));
y(5) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0));
y(4) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0))) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and b(2) and (not b(1)) and (not b(0)));
y(0) <= 
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and (not b(12)) and b(11) and b(10) and b(9) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and (not b(8)) and b(7) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and (not b(10)) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and b(7) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and (not b(13)) and b(12) and b(11) and b(10) and b(9) and (not b(8)) and b(7) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and (not b(10)) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and (not b(9)) and (not b(8)) and b(7) and b(6) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and (not b(11)) and b(10) and b(9) and b(8) and b(7) and b(6) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and (not b(9)) and (not b(8)) and b(7) and (not b(6)) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and (not b(12)) and b(11) and b(10) and b(9) and (not b(8)) and (not b(7)) and b(6) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and (not b(8)) and (not b(7)) and (not b(6)) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and (not b(9)) and b(8) and b(7) and b(6) and b(5) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and (not b(10)) and b(9) and b(8) and b(7) and (not b(6)) and b(5) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and (not b(9)) and b(8) and (not b(7)) and b(6) and b(5) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and (not b(11)) and b(10) and b(9) and b(8) and (not b(7)) and b(6) and (not b(5)) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and b(5) and b(4) and (not b(3)) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and (not b(10)) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and b(4) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and (not b(9)) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and b(3) and (not b(2)) and (not b(1)) and b(0)) or
		((not b(15)) and (not b(14)) and b(13) and b(12) and b(11) and b(10) and b(9) and b(8) and (not b(7)) and (not b(6)) and (not b(5)) and (not b(4)) and (not b(3)) and (not b(2)) and (not b(1)) and b(0));
END Behavioral;
